package as_pack;
    // Minimal RV64I parameter pack for templates
    parameter int reg_width = 64;
    parameter int instr_width = 32;
    parameter int imemdepth = 8192;
    parameter int dmemdepth = 1024;
    parameter int nr_gpios = 8;
    parameter int nr_regs = 32;
endpackage
