`timescale 1us/100ns

module tb;
    initial begin
        $dumpfile("../test.vcd");
        $dumpvars(0);
    end
endmodule
