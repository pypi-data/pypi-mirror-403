`timescale 1us/100ns

module tb;

endmodule
